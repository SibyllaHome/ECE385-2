module testRam (
					 input [7:0] read_addr,
					 input clk,
					 output logic [15:0] data_out);