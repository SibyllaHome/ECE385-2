module multiplier(input logic [7:0] SW,
						input logic [7:0] B,
						output logic [7:0] Aval
						output logic [7:0] Bval
						output logic X);

logic Q_, N;
logic [7:0] A,Q;

Q_ = 1'b0;	// Q_ initialize 0
Q  = B;		// Q  initialize to B
A  = 2'h00; // A  initialize 0000 0000 0000 0000

do
	begin
	if (Q[0] == 0 && Q_ == 0)
		begin
		
	
	
	
	
	
	end
while(N > 1'b0)				
						
						
						
						
						
						
endmodule
