module final_project_top_level(
										 
										 );
										 
										 
endmodule
