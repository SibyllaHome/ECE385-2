//------------------------------------------------------------------------------
// Company:          UIUC ECE Dept.
// Engineer:         Stephen Kempf
//
// Create Date:    17:44:03 10/08/06
// Design Name:    ECE 385 Lab 6 Given Code - Incomplete ISDU
// Module Name:    ISDU - Behavioral
//
// Comments:
//    Revised 03-22-2007
//    Spring 2007 Distribution
//    Revised 07-26-2013
//    Spring 2015 Distribution
//    Revised 02-13-2017
//    Spring 2017 Distribution
//------------------------------------------------------------------------------


module ISDU (   input logic         Clk, 
									Reset,
									Run,
									Continue,
									
				input logic[3:0]    Opcode, 
				input logic         IR_5,
				input logic         IR_11,
				input logic         BEN,
				  
				output logic        LD_MAR,
									LD_MDR,
									LD_IR,
									LD_BEN,
									LD_CC,
									LD_REG,
									LD_PC,
									LD_LED, // for PAUSE instruction
									
				output logic        GatePC,
									GateMDR,
									GateALU,
									GateMARMUX,
									
				output logic [1:0]  PCMUX,
				output logic        DRMUX,
									SR1MUX,
									SR2MUX,
									ADDR1MUX,
				output logic [1:0]  ADDR2MUX,
									ALUK,
				  
				output logic        Mem_CE,
									Mem_UB,
									Mem_LB,
									Mem_OE,
									Mem_WE
				);

	enum logic [4:0] {  Halted,
						LED_PAUSE1,LED_PAUSE2,
						S_18, 
						S_33_1, 
						S_33_2, 
						S_35, 
						S_32, 						// BEN
						S_01,							// ADD
						S_05,							// AND
						S_09, 						// NOT
						S_00, S_22, 				// BR
						S_12, 						// JMP
						S_04, S_21,					// JSR
						S_07,	S_23,	S_16_1, S_16_2, 		// STR
						S_06, S_25_1, S_25_2, S_27, Manual_Pause1, Manual_Pause2			// LDR
						}   State, Next_state;   // Internal state logic
		
	always_ff @ (posedge Clk)
	begin
		if (Reset) 
			State <= Halted;
		else 
			State <= Next_state;
	end
   
	always_comb
	begin 
		// Default next state is staying at current state
		Next_state = State;
		
		// Default controls signal values
		LD_MAR = 1'b0;
		LD_MDR = 1'b0;
		LD_IR = 1'b0;
		LD_BEN = 1'b0;
		LD_CC = 1'b0;
		LD_REG = 1'b0;
		LD_PC = 1'b0;
		LD_LED = 1'b0;
		 
		GatePC = 1'b0;
		GateMDR = 1'b0;
		GateALU = 1'b0;
		GateMARMUX = 1'b0;
		 
		ALUK = 2'b00;
		 
		PCMUX = 2'b00;
		DRMUX = 1'b0;
		SR1MUX = 1'b0;
		SR2MUX = 1'b0;
		ADDR1MUX = 1'b0;
		ADDR2MUX = 2'b00;
		 
		Mem_OE = 1'b1;
		Mem_WE = 1'b1;
	
		// Assign next state
		unique case (State)
			Halted : 
				if (Run) 
					Next_state = S_18;
					
//			Manual_Pause1:
//				if(~Continue)
//					Next_state = Manual_Pause1;
//				else
//					Next_state = Manual_Pause2;
//			Manual_Pause2:
//				if(Continue)
//					Next_state = Manual_Pause2;
//				else
//					Next_state = S_33_1;
					
			S_18 : 
				Next_state = S_33_1;

			// Any states involving SRAM require more than one clock cycles.
			// The exact number will be discussed in lecture.
			S_33_1 : 
				Next_state = S_33_2;
			S_33_2 : 
				Next_state = S_35;
			S_35 : 
				Next_state = S_32;

			S_32 : 									// BEN
				case (Opcode)
					4'b0001 : 						// ADD
						Next_state = S_01;
					4'b0101 :						// AND
						Next_state = S_05;
					4'b1001 :						// NOT
						Next_state = S_09;
					4'b0000 :						// BR
						Next_state = S_00;
					4'b1100 :						// JMP
						Next_state = S_12;
					4'b0100 :						// JSR
						Next_state = S_04;
					4'b0111 :						// STR
						Next_state = S_07;
					4'b0110 :						// LDR
						Next_state = S_06;		
					4'b1101 :						// Pause for LED
						Next_state = LED_PAUSE1;
						
						
					// You need to finish the rest of opcodes.....

					default : 
						Next_state = S_18;
				endcase
				
			S_01 : 
				Next_state = S_18;
			S_05 :
				Next_state = S_18;
			S_09 :
				Next_state = S_18;
			S_00 :
				if(BEN)
					Next_state = S_22; // can be 22 then to 18, or 18
				else
					Next_state = S_18;
			S_22 :
				Next_state = S_18;
			S_12 :
				Next_state = S_18;
			S_04 :
				Next_state = S_21; // can be 21, then to 18
			S_21 :
				Next_state = S_18;
			S_07 :
				Next_state = S_23; // 07 STR: MAR <- B + off6
			S_23 :
				Next_state = S_16_1; // 23 STR: MDR <- SR
			S_16_1:
				Next_state = S_16_2;
			S_16_2 :
				Next_state = S_18; // 16 STR: M[MAR] <- MDR
			S_06 :
				Next_state = S_25_1;
			S_25_1 :
				Next_state = S_25_2;
			S_25_2 :
				Next_state = S_27;
			S_27 :
				Next_state = S_18;
			
			// 2 LED PAUSE STATES
			LED_PAUSE1 :
				if(~Continue)
					Next_state = LED_PAUSE1;
				else
					Next_state = LED_PAUSE2;
			LED_PAUSE2 :
				if(Continue)
					Next_state = LED_PAUSE2;
				else
					Next_state = S_18;
			

			default : ;

		endcase
		
		// Assign control signals based on current state ///////////////////////////////////
		case (State)
		
		
			// SR1 MUX Select Bit : 0: IR[11:9]
			//                      1: IR[8 :6]
			
			// DR MUX Select Bit :	0: IR[11:9]
			//								1: 3'b111
			
			// SR2 MUX Select Bit:	0: SR2_OUT
			//								1: 5-bits SEXT
		
		
		
			Halted: ;	// do nothing
			
			S_18 :  //MAR<-PC; PC<-PC+1
				begin 
					GatePC = 1'b1;
					LD_MAR = 1'b1;
					PCMUX = 2'b10;
					LD_PC = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end

			S_33_1 : //MDR<-M(MAR)
				begin
					Mem_OE = 1'b0;
					Mem_WE = 1'b1;
				end
				
			S_33_2 : //MDR<-M(MAR)
				begin 
					Mem_OE = 1'b0;
					Mem_WE = 1'b1;
					
					LD_MDR = 1'b1;
				end
				
			S_35 : //IR<-MDR
				begin 
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
					
					GateMDR = 1'b1;
					LD_IR = 1'b1;
				end
				
			S_32 : //BEN
				LD_BEN = 1'b1;
				
			S_01 : //ADD
				begin 
					SR2MUX = IR_5; 
					SR1MUX = 1'b1;
					ALUK = 2'b00;
					GateALU = 1'b1;
					LD_REG = 1'b1;
					LD_CC = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_05 : //AND DR<-SR1 & OP2, set CC
				begin
					SR2MUX = IR_5;
					SR1MUX = 1'b1;
					ALUK = 2'b01;
					GateALU = 1'b1;
					LD_REG = 1'b1;
					LD_CC = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_09 :	//NOT DR<-NOT(SR), set CC
				begin
					SR1MUX = 1'b1;
					ALUK = 2'b10;
					GateALU = 1'b1;
					LD_REG = 1'b1;
					LD_CC = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_00 : //BEN
				begin
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_22 : //PC<-PC+off9
				begin
					ADDR2MUX = 2'b01; //IR[8:0]
					ADDR1MUX = 1'b1;	//PC
					PCMUX = 2'b01;   //add
					LD_PC = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_12 : //PC<-BaseR
				begin
					SR1MUX = 1'b1;
					LD_PC = 1'b1;
					PCMUX = 2'b01;
					ADDR1MUX = 1'b0;
					ADDR2MUX = 2'b11;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_04 : //R7<-PC
				begin
					GatePC = 1'b1;
					DRMUX = IR_11;
					LD_REG = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_21 : //PC<-PC+off11
				begin
					LD_PC = 1'b1;
					ADDR2MUX = 2'b00;
					ADDR1MUX = 1'b1; //PC
					PCMUX = 2'b01;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_07 : //MAR<-B+off6
				begin
					SR1MUX = 1'b1;
					ADDR1MUX = 1'b0;
					ADDR2MUX = 2'b10;
					GateMARMUX = 1'b1;
					LD_MAR = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_23 : // MDR<-SR
				begin
					SR1MUX = 1'b0;
					ALUK = 2'b11; // pass
					GateALU = 1'b1;
					LD_MDR = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_16_1 : // M[MAR]<-MDR
				begin
					Mem_OE = 1'b1;
					Mem_WE = 1'b0;
				end
				
			S_16_2 :
				begin
					Mem_OE = 1'b1;
					Mem_WE = 1'b0;
				end
				
			S_06 : // MAR<-B+off6
				begin
					SR1MUX = 1'b1;
					ADDR1MUX = 1'b0;
					ADDR2MUX = 2'b10;
					GateMARMUX = 1'b1;
					LD_MAR = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			S_25_1: //MDR<-M[MAR]
				begin
					Mem_OE = 1'b0;
					Mem_WE = 1'b1;
				end
				
			S_25_2 :
				begin
					Mem_OE = 1'b0;
					Mem_WE = 1'b1;
					LD_MDR = 1'b1;
				end
				
			S_27: //DR<-MDR, set CC
				begin
					DRMUX = 1'b0;
					LD_REG = 1'b1;
					LD_CC = 1'b1;
					GateMDR = 1'b1;
					
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			LED_PAUSE1:
				begin
					LD_LED = 1'b1;
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end
				
			LED_PAUSE2:
				begin
					Mem_OE = 1'b1;
					Mem_WE = 1'b1;
				end

				
			default :
			begin
				Mem_OE = 1'b1;
				Mem_WE = 1'b1;
			end
			
		endcase
	end 

		// always active
	assign Mem_CE = 1'b0;
	assign Mem_UB = 1'b0;
	assign Mem_LB = 1'b0;
	
endmodule
